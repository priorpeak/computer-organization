`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/09/2021 09:59:39 PM
// Design Name: 
// Module Name: mov1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mov1(out, in);
    // Input (Source register)
    input  in;
    
    // Output (Destination register)
    output out;
    
    assign out = in;
endmodule
